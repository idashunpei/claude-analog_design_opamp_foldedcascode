* Folded Cascode OTA — Transient (Unity-Gain Feedback)
.model nch nmos level=1 vto=0.5 kp=0.0002
+ lambda=0.1
.model pch pmos level=1 vto=-0.5 kp=8e-05
+ lambda=0.15

* --- Supply & Bias ---
VDD   vdd   0   1.8
Vbias vbias 0   1.1000
Vcn   vcn   0   1.3000
Vbp   vbp   0   1.1000
Vcp   vcp   0   0.9000

* --- Step input on non-inverting input ---
Vinp  vinp  0  PULSE(0.5 1.3 0.5u 1n 1n 4u 8u)
* --- OTA core (vinn = vout for unity-gain feedback) ---
M0   vtail  vbias  vdd  vdd  pch  W=31.25u  L=0.50u
M1   na     vinp   vtail vdd pch  W=24.67u  L=0.50u
M2   vout   vout   vtail vdd pch  W=24.67u  L=0.50u
M3   na     vcn    nc    0   nch  W=22.22u  L=0.50u
M4   vout   vcn    nd    0   nch  W=22.22u  L=0.50u
M5   nc     nc     0     0   nch  W=22.22u  L=0.50u
M6   nd     nc     0     0   nch  W=22.22u  L=0.50u
M7   na     vcp    ne    vdd pch  W=15.62u  L=0.50u
M8   vout   vcp    nf    vdd pch  W=15.62u  L=0.50u
M9   ne     vbp    vdd   vdd pch  W=15.62u  L=0.50u
M10  nf     vbp    vdd   vdd pch  W=15.62u L=0.50u
CL   vout   0      2e-12
.control
    tran 1n 10u
    wrdata tran_fb_out v(vout) v(vinp)
    quit
.endc
.end
