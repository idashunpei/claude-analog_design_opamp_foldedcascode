* Folded Cascode OTA — AC Analysis
.model nch nmos level=1 vto=0.5 kp=0.0002
+ lambda=0.1
.model pch pmos level=1 vto=-0.5 kp=8e-05
+ lambda=0.15

* --- Supply & Bias ---
VDD   vdd   0   1.8
Vbias vbias 0   1.1000
Vbn   vbn   0   0.7000
Vcn   vcn   0   0.9000
Vbp   vbp   0   1.1000
Vcp   vcp   0   0.9000

* --- Differential AC input ---
Vinp  vinp  0  DC 0.9  AC  0.5
Vinn  vinn  0  DC 0.9  AC -0.5
* --- OTA core ---
M0   vtail  vbias  vdd  vdd  pch  W=31.25u  L=0.50u
M1   na     vinp   vtail vdd pch  W=24.67u  L=0.50u
M2   vout   vinn   vtail vdd pch  W=24.67u  L=0.50u
M3   na     vcn    nc    0   nch  W=12.50u  L=0.50u
M4   vout   vcn    nd    0   nch  W=12.50u  L=0.50u
M5   nc     vbn    0     0   nch  W=12.50u  L=0.50u
M6   nd     vbn    0     0   nch  W=12.50u  L=0.50u
M7   na     vcp    ne    vdd pch  W=15.62u  L=0.50u
M8   vout   vcp    nf    vdd pch  W=15.62u  L=0.50u
M9   ne     vbp    vdd   vdd pch  W=15.62u  L=0.50u
M10  nf     vbp    vdd   vdd pch  W=15.62u L=0.50u
* --- Load ---
CL   vout   0      2e-12

* --- DC-feedback inductor: short at DC, open at AC ---
Lfb   vout  vinn  1T
.control
    ac dec 100 1 10G
    wrdata ac_out v(vout)
    quit
.endc
.end
